LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY banco_de_registradores_tb IS
END ENTITY;

ARCHITECTURE a_banco_de_registradores_tb OF banco_de_registradores_tb IS
    COMPONENT banco_de_registradores
    END ARCHITECTURE;